CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 84 1918 1006
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 180 457 277
42991634 0
0
6 Title:
5 Name:
0
0
0
31
4 4511
219 824 286 0 1 29
0 0
0
0 0 4832 0
4 4511
-14 -60 14 -52
2 U6
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 0 0 0 0
1 U
5130 0 0
2
45439.3 0
0
13 Logic Switch~
5 251 779 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 253 700 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90125e-315 5.32571e-315
0
13 Logic Switch~
5 254 737 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90125e-315 5.30499e-315
0
13 Logic Switch~
5 250 624 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90125e-315 5.26354e-315
0
13 Logic Switch~
5 252 660 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 241 459 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90125e-315 5.32571e-315
0
13 Logic Switch~
5 245 572 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90125e-315 5.30499e-315
0
13 Logic Switch~
5 244 535 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90125e-315 5.26354e-315
0
13 Logic Switch~
5 243 495 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 240 288 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90125e-315 5.30499e-315
0
13 Logic Switch~
5 242 324 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90125e-315 5.26354e-315
0
13 Logic Switch~
5 244 401 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 243 364 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 325 117 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
5.90125e-315 5.32571e-315
0
13 Logic Switch~
5 327 153 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3670 0 0
2
5.90125e-315 5.30499e-315
0
13 Logic Switch~
5 329 230 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5616 0 0
2
5.90125e-315 5.26354e-315
0
13 Logic Switch~
5 328 193 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9323 0 0
2
5.90125e-315 0
0
7 Ground~
168 1022 119 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
317 0 0
2
45439.3 0
0
9 CA 7-Seg~
184 1120 188 0 18 19
10 37 38 39 40 41 42 43 44 45
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
6 BLUECA
13 -41 55 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3108 0 0
2
45439.3 0
0
9 CC 7-Seg~
183 1022 162 0 13 19
10 11 10 9 12 8 7 6 5 2
1 1 1 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
4299 0 0
2
5.90125e-315 0
0
5 4030~
219 400 732 0 3 22
0 29 3 25
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
9672 0 0
2
5.90125e-315 5.32571e-315
0
5 4030~
219 398 693 0 3 22
0 30 3 26
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7876 0 0
2
5.90125e-315 0
0
5 4030~
219 399 646 0 3 22
0 31 3 27
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
6369 0 0
2
5.90125e-315 0
0
5 4030~
219 400 597 0 3 22
0 32 3 28
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
9172 0 0
2
5.90125e-315 0
0
5 4030~
219 401 561 0 3 22
0 33 3 13
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
7100 0 0
2
5.90125e-315 0
0
5 4030~
219 398 521 0 3 22
0 34 3 14
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3820 0 0
2
5.90125e-315 0
0
5 4030~
219 399 481 0 3 22
0 35 3 15
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
7678 0 0
2
5.90125e-315 0
0
5 4030~
219 399 440 0 3 22
0 36 3 16
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
961 0 0
2
5.90125e-315 0
0
6 74LS83
105 603 503 0 14 29
0 24 23 22 21 28 27 26 25 4
8 7 6 5 46
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3178 0 0
2
5.90125e-315 0
0
6 74LS83
105 656 222 0 14 29
0 20 19 18 17 16 15 14 13 3
11 10 9 12 4
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3409 0 0
2
5.90125e-315 0
0
39
2 0 3 0 0 4096 0 22 0 0 31 2
384 741
334 741
1 0 3 0 0 4096 0 2 0 0 31 2
263 779
336 779
14 9 4 0 0 8320 0 31 30 0 0 5
688 267
701 267
701 574
571 574
571 548
1 9 2 0 0 4224 0 19 21 0 0 2
1022 127
1022 120
13 8 5 0 0 4224 0 30 21 0 0 3
635 521
1043 521
1043 198
12 7 6 0 0 4224 0 30 21 0 0 3
635 512
1037 512
1037 198
11 6 7 0 0 4224 0 30 21 0 0 3
635 503
1031 503
1031 198
10 5 8 0 0 4224 0 30 21 0 0 3
635 494
1025 494
1025 198
3 8 13 0 0 8320 0 26 31 0 0 4
434 561
441 561
441 249
624 249
3 7 14 0 0 8320 0 27 31 0 0 4
431 521
458 521
458 240
624 240
3 6 15 0 0 8320 0 28 31 0 0 6
432 481
468 481
468 237
563 237
563 231
624 231
3 5 16 0 0 8320 0 29 31 0 0 4
432 440
448 440
448 222
624 222
1 4 17 0 0 4224 0 17 31 0 0 4
341 230
548 230
548 213
624 213
1 3 18 0 0 4224 0 18 31 0 0 4
340 193
560 193
560 204
624 204
1 2 19 0 0 4224 0 16 31 0 0 4
339 153
579 153
579 195
624 195
1 1 20 0 0 4224 0 15 31 0 0 4
337 117
591 117
591 186
624 186
1 4 21 0 0 4224 0 13 30 0 0 4
256 401
501 401
501 494
571 494
1 3 22 0 0 4224 0 14 30 0 0 4
255 364
520 364
520 485
571 485
1 2 23 0 0 4224 0 12 30 0 0 4
254 324
531 324
531 476
571 476
1 1 24 0 0 4224 0 11 30 0 0 4
252 288
546 288
546 467
571 467
3 8 25 0 0 8320 0 22 30 0 0 4
433 732
513 732
513 530
571 530
3 7 26 0 0 8320 0 23 30 0 0 4
431 693
495 693
495 521
571 521
3 6 27 0 0 8320 0 24 30 0 0 4
432 646
480 646
480 512
571 512
3 5 28 0 0 12416 0 25 30 0 0 4
433 597
470 597
470 503
571 503
0 2 3 0 0 0 0 0 29 26 0 3
334 490
334 449
383 449
0 2 3 0 0 0 0 0 28 27 0 3
334 530
334 490
383 490
0 2 3 0 0 0 0 0 27 28 0 3
334 569
334 530
382 530
0 2 3 0 0 0 0 0 26 29 0 4
334 606
334 569
385 569
385 570
0 2 3 0 0 0 0 0 25 30 0 3
334 657
334 606
384 606
0 2 3 0 0 0 0 0 24 31 0 3
334 704
334 655
383 655
9 2 3 0 0 12416 0 31 23 0 0 7
624 267
624 292
731 292
731 779
334 779
334 702
382 702
1 1 29 0 0 12416 0 4 22 0 0 4
266 737
274 737
274 723
384 723
1 1 30 0 0 12416 0 3 23 0 0 4
265 700
277 700
277 684
382 684
1 1 31 0 0 12416 0 6 24 0 0 4
264 660
277 660
277 637
383 637
1 1 32 0 0 12416 0 5 25 0 0 4
262 624
278 624
278 588
384 588
1 1 33 0 0 12416 0 8 26 0 0 4
257 572
269 572
269 552
385 552
1 1 34 0 0 12416 0 9 27 0 0 4
256 535
273 535
273 512
382 512
1 1 35 0 0 12416 0 10 28 0 0 4
255 495
278 495
278 472
383 472
1 1 36 0 0 12416 0 7 29 0 0 4
253 459
282 459
282 431
383 431
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
187 390 232 414
197 398 221 414
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
187 243 232 267
197 251 221 267
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
276 220 321 244
286 228 310 244
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
277 77 322 101
287 85 311 101
3 MSB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
